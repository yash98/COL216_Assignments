library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
library UNISIM;  

entity Actrl is
    port (
        ins27_21: in std_logic_vector(7 downto 0);
        --op: out std_logic_vector();
    );    
end entity;